module(SDCLK, Reset);
	
endmodule;