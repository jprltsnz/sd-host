   module remap(
                    input logic [2047:0] mem_data_out,
                    output logic [15:0]  sdma_address_low,
                    output logic [15:0]  sdma_address_high,
                    output logic [15:0]  block_size,
                    output logic [15:0]  block_count,
                    output logic [15:0]  argument_0,
                    output logic [15:0]  argument_1,
                    output logic [15:0]  response_0,
                    output logic [15:0]  response_1,
                    output logic [15:0]  response_2,
                    output logic [15:0]  response_3,
                    output logic [15:0]  response_4,
                    output logic [15:0]  response_5,
                    output logic [15:0]  response_6,
                    output logic [15:0]  response_7,
                    output logic [15:0]  buffer_data_port_0,
                    output logic [15:0]  buffer_data_port_1,
                    output logic [31:0]  present_state,
                    output logic [7:0]   host_control,
                    output logic [7:0]   power_control,
                    output logic [7:0]   block_gap_control,
                    output logic [7:0]   wakeup_control,
                    output logic [15:0]  clock_control,
                    output logic [7:0]   timeout_control,
                    output logic [7:0]   software_reset,
                    output logic [15:0]  normal_interrupt_status,
                    output logic [15:0]  error_interruprt_status,
                    output logic [15:0]  normal_interrupt_status_en,
                    output logic [15:0]  error_interruprt_status_en,
                    output logic [15:0]  normal_interrupt_signal_en,
                    output logic [15:0]  error_interruprt_signal_en,
                    output logic [15:0]  auto_cmd_12_error_status,
                    output logic [31:0]  capabilities,
                    output logic [15:0]  capabilities_resrv,
                    output logic [31:0]  max_current_capabilities,
                    output logic [31:0]  max_current_capabilities_resrv,
                    output logic [15:0]  force_event_auto_cmd_12_error_status,
                    output logic [15:0]  force_event_error_interrupt_status,
                    output logic [8:0]   adma_error_status,
                    output logic [63:0]  adma_system_address,
                    output logic [15:0]  slot_interrupt_status,
                    output logic [15:0]  host_controller_version
                    );

   assign sdma_address_low = mem_data_out[15:0];
   assign sdma_address_high = mem_data_out[31:16];
   assign block_size = mem_data_out[47:32];
   assign block_count = mem_data_out[63:48];
   assign argument_0 = mem_data_out[79:64];
   assign argument_1 = mem_data_out[95:80];
   assign response_0 = mem_data_out[111:96];
   assign response_1 = mem_data_out[127:112];
   assign response_2 = mem_data_out[143:128];
   assign response_3 = mem_data_out[159:144];
   assign response_4 = mem_data_out[175:160];
   assign response_5 = mem_data_out[191:176];
   assign response_6 = mem_data_out[207:192];
   assign response_7 = mem_data_out[223:208];
   assign buffer_data_port_0 = mem_data_out[239:224];
   assign buffer_data_port_1 = mem_data_out[255:240];
   assign present_state = mem_data_out[271:256];
   assign host_control = mem_data_out[287:272];
   assign power_control = mem_data_out[303:288];
   assign block_gap_control = mem_data_out[319:304];
   assign wakeup_control = mem_data_out[335:320];
   assign clock_control = mem_data_out[351:336];
   assign timeout_control = mem_data_out[367:352];
   assign software_reset = mem_data_out[383:368];
   assign normal_interrupt_status = mem_data_out[399:384];
   assign error_interruprt_status = mem_data_out[415:400];
   assign normal_interrupt_status_en = mem_data_out[431:416];
   assign error_interruprt_status_en = mem_data_out[447:432];
   assign normal_interrupt_signal_en = mem_data_out[463:448];
   assign error_interruprt_signal_en = mem_data_out[479:464];
   assign auto_cmd_12_error_status = mem_data_out[495:480];
   assign capabilities = mem_data_out[543:512];
   assign capabilities_resrv = mem_data_out[575:544];
   assign max_current_capabilities = mem_data_out[607:576];
   assign max_current_capabilities_resrv = mem_data_out[639:608];
   assign force_event_auto_cmd_12_error_status = mem_data_out[655:640];
   assign force_event_error_interrupt_status = mem_data_out[671:656];
   assign adma_error_status = mem_data_out[679:672];
   assign adma_system_address = mem_data_out[767:704];
   assign slot_interrupt_status = mem_data_out[2031:2016];
   assign host_controller_version = mem_data_out[2047:2032];
endmodule // remap
