module(reset, in, out, new_set);
	
	parameter BITS = 48;
	
	input wire reset, in, new_set;
	output wire [BITS-1:0] out;
	
	
endmodule